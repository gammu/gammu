Gammu All Mobile Management Utilities - Installation
====================================================

Se docs/manual/project/install.rst för installationsguiden eller se kapitlet ”Kompilera Gammu” i Gammu-manualen.
