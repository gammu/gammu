Gammu All Mobile Management Utilities (Gammu alla mobilhanteringsverktyg)
=========================================================================

Gammu är ett bibliotek och kommandoradsverktyg för mobiltelefoner. Det
publiceras under GNU GPL version 2.

Det påbörjades av Marcin Wiacek och andra. Från början baserades koden på
Gnokii <https://www.gnokii.org/>- och senare MyGnokii
<http://www.mwiacek.com/>-projekten. Gammu kallades (fram till version 0.58)
för MyGnokii2.

För närvarande är leds projektet av Michael Cihar <michal@cihar.com> med
hjälp från många bidragsgivare.

.. bild:: https://travis-ci.org/gammu/gammu.svg?branch=master
    :alt: Byggstatus :target: https://travis-ci.org/gammu/gammu

.. bild:: https://ci.appveyor.com/api/projects/status/dkm2eam66rbhhuwn/branch/master?svg=true
    :alt: Byggstatus för Windows :target:
    https://ci.appveyor.com/project/nijel/gammu/branch/master

.. bild:: https://hosted.weblate.org/widgets/gammu/-/svg-badge.svg
    :alt: Översättningsstatus :target:
    https://hosted.weblate.org/engage/gammu/?utm_source=widget

.. bild:: https://scan.coverity.com/projects/2890/badge.svg?flat=1
    :alt: Coverity-genomsökning :target: https://scan.coverity.com/projects/2890

.. bild:: https://img.shields.io/liberapay/receives/Gammu.svg
    :alt: Liberapay :target: https://liberapay.com/Gammu/donate

.. bild:: https://www.bountysource.com/badge/team?team_id=23177&style=bounties_received
    :alt: Bountysource :target:
    https://www.bountysource.com/teams/gammu/issues?utm_source=Gammu&utm_medium=shield&utm_campaign=bounties_received

Vidare information
==================

Du kan hitta vidare information på <https://wammu.eu/gammu/>.

Det finns också en Gammu-manual tillgänglig i docs/manual. Du kan bygga
HTML-versionen av den med hjälp av make manual-html vilken också går att
läsa på <https://wammu.eu/docs/manual/>.


Återkoppling och felrapporter
=============================

All möjlig återkoppling är välkommen, se <https://wammu.eu/support/> för
information om hur du kontaktar utvecklarna.


Stöd utvecklarna
================

Du kan ge uppskattning till utvecklarna via <https://wammu.eu/donate/>.
